module decoder()


endmodule
